.param Tox = 1e-09

.param Toxe1 = 'Tox + 2.5e-10' $ 1.25e-09
.param Toxp1 = 'Tox' $ 1e-09
.param Toxm1 = 'Toxe1' $ 1.25e-09
.param dTox1 = 'Toxe1 - Toxp1' $ 2.5e-10
.param Toxref1 = 'Toxe1' $ 1.25e-09

.param Toxe2 = 'Tox + 3e-10' $ 1.3e-09
.param Toxp2 = 'Tox' $ 1e-09
.param Toxm2 = 'Toxe2' $ 1.3e-09
.param dTox2 = 'Toxe2 - Toxp2' $ 3e-10
.param Toxref2 = 'Toxe2' $ 1.3e-09

.model nmos nmos
+ a0 = 1
+ a1 = 0
+ a2 = 1
+ acde = 1
+ acnqsmod = 0
+ agidl = 0.0002
+ ags = 0
+ aigbacc = 0.012
+ aigbinv = 0.014
+ aigc = 0.02
+ aigsd = 0.02
+ alpha0 = 0.074
+ alpha1 = 0.005
+ at = 33000
+ b0 = 0
+ b1 = 0
+ beta0 = 30
+ bgidl = 2.1e+09
+ bigbacc = 0.0028
+ bigbinv = 0.004
+ bigc = 0.0025
+ bigsd = 0.0025
+ binunit = 1
+ bvd = 10
+ bvs = 10
+ capmod = 2
+ cdsc = 0
+ cdscb = 0
+ cdscd = 0
+ cgbo = 2.56e-11
+ cgdl = 2.653e-10
+ cgdo = 1.1e-10
+ cgidl = 0.0002
+ cgsl = 2.653e-10
+ cgso = 1.1e-10
+ cigbacc = 0.002
+ cigbinv = 0.004
+ cigc = 0.002
+ cigsd = 0.002
+ cit = 0
+ cjd = 0.0005
+ cjs = 0.0005
+ cjswd = 5e-10
+ cjswgd = 5e-10
+ cjswgs = 3e-10
+ cjsws = 5e-10
+ ckappad = 0.03
+ ckappas = 0.03
+ delta = 0.01
+ diomod = 1
+ dmcg = 0
+ dmcgt = 0
+ dmci = 0
+ dmdg = 0
+ drout = 0.5
+ dsub = 0.1
+ dtox = 'dTox1'
+ dvt0 = 1
+ dvt0w = 0
+ dvt1 = 2
+ dvt1w = 0
+ dvt2 = 0
+ dvt2w = 0
+ dvtp0 = 1e-10
+ dvtp1 = 0.1
+ dwb = 0
+ dwg = 0
+ dwj = 0
+ egidl = 0.8
+ eigbinv = 1.1
+ epsrox = 3.9
+ eta0 = 0.0055
+ etab = 0
+ fnoimod = 1
+ fprout = 0.2
+ gbmin = 1e-10
+ geomod = 1
+ igbmod = 1
+ igcmod = 1
+ ijthdfwd = 0.01
+ ijthdrev = 0.001
+ ijthsfwd = 0.01
+ ijthsrev = 0.001
+ jsd = 0.0001
+ jss = 0.0001
+ jswd = 1e-11
+ jswgd = 1e-10
+ jswgs = 1e-10
+ jsws = 1e-11
+ k1 = 0.4
+ k2 = 0
+ k3 = 0
+ k3b = 0
+ keta = 0.04
+ kt1 = -0.11
+ kt1l = 0
+ kt2 = 0.022
+ level = 54
+ lint = 3.75e-09
+ ll = 0
+ lln = 1
+ lpe0 = 0
+ lpeb = 0
+ lw = 0
+ lwl = 0
+ lwn = 1
+ minv = 0.05
+ mjd = 0.5
+ mjs = 0.5
+ mjswd = 0.33
+ mjswgd = 0.33
+ mjswgs = 0.33
+ mjsws = 0.33
+ mobmod = 0
+ moin = 15
+ ndep = 3.24e+18
+ nfactor = 2.22
+ ngate = 1e+23
+ ngcon = 1
+ nigbacc = 1
+ nigbinv = 3
+ nigc = 1
+ njd = 1
+ njs = 1
+ noff = 0.9
+ nsd = 2e+20
+ ntox = 1
+ paramchk = 1
+ pbd = 1
+ pbs = 1
+ pbswd = 1
+ pbswgd = 1
+ pbswgs = 1
+ pbsws = 1
+ pclm = 0.02
+ pdiblc1 = 0.001
+ pdiblc2 = 0.001
+ pdiblcb = -0.005
+ pdits = 0.08
+ pditsd = 0.23
+ pditsl = 2.3e+06
+ permod = 1
+ phin = 0
+ pigcd = 1
+ poxedge = 1
+ prt = 0
+ prwb = 0
+ prwg = 0
+ pscbe1 = 8.14e+08
+ pscbe2 = 1e-07
+ pvag = 1e-20
+ rbdb = 15
+ rbodymod = 1
+ rbpb = 5
+ rbpd = 15
+ rbps = 15
+ rbsb = 15
+ rdsmod = 0
+ rdsw = 155
+ rdswmin = 0
+ rdw = 80
+ rdwmin = 0
+ rgatemod = 1
+ rsh = 5
+ rshg = 0.4
+ rsw = 80
+ rswmin = 0
+ tcj = 0.001
+ tcjsw = 0.001
+ tcjswg = 0.001
+ tnoimod = 0
+ tnom = 27
+ toxe = 'Toxe1'
+ toxm = 'Toxm1'
+ toxp = 'Toxp1'
+ toxref = 'Toxref1'
+ tpb = 0.005
+ tpbsw = 0.005
+ tpbswg = 0.005
+ trnqsmod = 0
+ u0 = 0.054
+ ua = 6e-10
+ ua1 = 4.31e-09
+ ub = 1.2e-18
+ ub1 = 7.61e-18
+ uc = 0
+ uc1 = -5.6e-11
+ ute = -1.5
+ version = 4
+ vfb = -0.55
+ voff = -0.13
+ voffcv = 0.02
+ voffl = 0
+ vsat = 170000
+ vth0 = 0.46893
+ w0 = 2.5e-06
+ wint = 5e-09
+ wl = 0
+ wln = 1
+ wr = 1
+ ww = 0
+ wwl = 0
+ wwn = 1
+ xgl = 0
+ xgw = 0
+ xj = 1.4e-08
+ xjbvd = 1
+ xjbvs = 1
+ xl = -2e-08
+ xpart = 0
+ xrcrg1 = 12
+ xrcrg2 = 5
+ xtid = 3
+ xtis = 3

.model pmos pmos
+ a0 = 1
+ a1 = 0
+ a2 = 1
+ acde = 1
+ acnqsmod = 0
+ agidl = 0.0002
+ ags = 1e-20
+ aigbacc = 0.012
+ aigbinv = 0.014
+ aigc = 0.010687
+ aigsd = 0.010687
+ alpha0 = 0.074
+ alpha1 = 0.005
+ at = 33000
+ b0 = 0
+ b1 = 0
+ beta0 = 30
+ bgidl = 2.1e+09
+ bigbacc = 0.0028
+ bigbinv = 0.004
+ bigc = 0.0012607
+ bigsd = 0.0012607
+ binunit = 1
+ bvd = 10
+ bvs = 10
+ capmod = 2
+ cdsc = 0
+ cdscb = 0
+ cdscd = 0
+ cgbo = 2.56e-11
+ cgdl = 2.653e-10
+ cgdo = 1.1e-10
+ cgidl = 0.0002
+ cgsl = 2.653e-10
+ cgso = 1.1e-10
+ cigbacc = 0.002
+ cigbinv = 0.004
+ cigc = 0.0008
+ cigsd = 0.0008
+ cit = 0
+ cjd = 0.0005
+ cjs = 0.0005
+ cjswd = 5e-10
+ cjswgd = 5e-10
+ cjswgs = 3e-10
+ cjsws = 5e-10
+ ckappad = 0.03
+ ckappas = 0.03
+ delta = 0.01
+ diomod = 1
+ dmcg = 0
+ dmcgt = 0
+ dmci = 0
+ dmdg = 0
+ drout = 0.56
+ dsub = 0.1
+ dtox = 'dTox2'
+ dvt0 = 1
+ dvt0w = 0
+ dvt1 = 2
+ dvt1w = 0
+ dvt2 = -0.032
+ dvt2w = 0
+ dvtp0 = 1e-11
+ dvtp1 = 0.05
+ dwb = 0
+ dwg = 0
+ dwj = 0
+ egidl = 0.8
+ eigbinv = 1.1
+ epsrox = 3.9
+ eta0 = 0.0055
+ etab = 0
+ fnoimod = 1
+ fprout = 0.2
+ gbmin = 1e-10
+ geomod = 1
+ igbmod = 1
+ igcmod = 1
+ ijthdfwd = 0.01
+ ijthdrev = 0.001
+ ijthsfwd = 0.01
+ ijthsrev = 0.001
+ jsd = 0.0001
+ jss = 0.0001
+ jswd = 1e-11
+ jswgd = 1e-10
+ jswgs = 1e-10
+ jsws = 1e-11
+ k1 = 0.4
+ k2 = -0.01
+ k3 = 0
+ k3b = 0
+ keta = -0.047
+ kt1 = -0.11
+ kt1l = 0
+ kt2 = 0.022
+ level = 54
+ lint = 3.75e-09
+ ll = 0
+ lln = 1
+ lpe0 = 0
+ lpeb = 0
+ lw = 0
+ lwl = 0
+ lwn = 1
+ minv = 0.05
+ mjd = 0.5
+ mjs = 0.5
+ mjswd = 0.33
+ mjswgd = 0.33
+ mjswgs = 0.33
+ mjsws = 0.33
+ mobmod = 0
+ moin = 15
+ ndep = 2.44e+18
+ nfactor = 2.1
+ ngate = 1e+23
+ ngcon = 1
+ nigbacc = 1
+ nigbinv = 3
+ nigc = 1
+ njd = 1
+ njs = 1
+ noff = 0.9
+ nsd = 2e+20
+ ntox = 1
+ paramchk = 1
+ pbd = 1
+ pbs = 1
+ pbswd = 1
+ pbswgd = 1
+ pbswgs = 1
+ pbsws = 1
+ pclm = 0.12
+ pdiblc1 = 0.001
+ pdiblc2 = 0.001
+ pdiblcb = 3.4e-08
+ pdits = 0.08
+ pditsd = 0.23
+ pditsl = 2.3e+06
+ permod = 1
+ phin = 0
+ pigcd = 1
+ poxedge = 1
+ prt = 0
+ prwb = 0
+ prwg = 0
+ pscbe1 = 8.14e+08
+ pscbe2 = 9.58e-07
+ pvag = 1e-20
+ rbdb = 15
+ rbodymod = 1
+ rbpb = 5
+ rbpd = 15
+ rbps = 15
+ rbsb = 15
+ rdsmod = 0
+ rdsw = 155
+ rdswmin = 0
+ rdw = 75
+ rdwmin = 0
+ rgatemod = 1
+ rsh = 5
+ rshg = 0.4
+ rsw = 75
+ rswmin = 0
+ tcj = 0.001
+ tcjsw = 0.001
+ tcjswg = 0.001
+ tnoimod = 0
+ tnom = 27
+ toxe = 'Toxe2'
+ toxm = 'Toxm2'
+ toxp = 'Toxp2'
+ toxref = 'Toxref2'
+ tpb = 0.005
+ tpbsw = 0.005
+ tpbswg = 0.005
+ trnqsmod = 0
+ u0 = 0.02
+ ua = 2e-09
+ ua1 = 4.31e-09
+ ub = 5e-19
+ ub1 = 7.61e-18
+ uc = 0
+ uc1 = -5.6e-11
+ ute = -1.5
+ version = 4
+ vfb = 0.55
+ voff = -0.126
+ voffcv = 0.02
+ voffl = 0
+ vsat = 150000
+ vth0 = -0.49158
+ w0 = 2.5e-06
+ wint = 5e-09
+ wl = 0
+ wln = 1
+ wr = 1
+ ww = 0
+ wwl = 0
+ wwn = 1
+ xgl = 0
+ xgw = 0
+ xj = 1.4e-08
+ xjbvd = 1
+ xjbvs = 1
+ xl = -2e-08
+ xpart = 0
+ xrcrg1 = 12
+ xrcrg2 = 5
+ xtid = 3
+ xtis = 3

