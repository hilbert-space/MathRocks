.param L = 50n

.param Tox = 1n

.param nToxe   = 'Tox + 0.63n'   $ 1.63
.param nToxp   = 'Tox'           $ 1n
.param nToxm   = 'nToxe'         $ 1.63
.param nToxref = 'nToxe'         $ 1.63
.param ndTox   = 'nToxe - nToxp' $ 0.63n

.param pToxe   = 'Tox + 0.6n'    $ 1.6n
.param pToxp   = 'Tox'           $ 1n
.param pToxm   = 'pToxe'         $ 1.6n
.param pToxref = 'pToxe'         $ 1.6n
.param pdTox   = 'pToxe - pToxp' $ 0.6n

* INV_X1

* Generated by: xspice 3.06 28-Mar-2013
* Date: 29-Sep-2013 16:09:04
* Path: /home/ivauk/Research/SPACE/inverter
* Language: SPICE

.subckt INV_X1 pbulk nbulk A VDD VSS ZN
m1 ZN A VSS SUBSTR NMOS_VTH w=90n l='L' ad=9.45f pd=300n nrd=1.1667 as=9.45f
+  ps=300n nrs=1.1667
m2 ZN A VDD 1 PMOS_VTH w=135n l='L' ad=14.175f pd=345n nrd=777.78m as=14.175f
+  ps=345n nrs=777.78m
.ends INV_X1

.model NMOS_VTH nmos level=54 tnom=27 epsrox=3.9 eta0=8m nfactor=1.6 wint=5n
+  cgso=110p cgdo=110p toxe='nToxe' toxp='nToxp' toxm='nToxm' toxref='nToxref' dtox='ndTox'
+  lint=3.75n vth0=607.8m k1=400m u0=50m vsat=170k rdsw=155 ndep=3.24e18
+  xj=19.8n version=4.0 binunit=1 paramchk=1 mobmod=0 capmod=2 igcmod=1
+  igbmod=1 geomod=1 diomod=1 rdsmod=0 rbodymod=1 rgatemod=1 permod=1
+  acnqsmod=0 trnqsmod=0 ll=0 wl=0 lln=1 wln=1 lw=0 ww=0 lwn=1 wwn=1 lwl=0
+  wwl=0 xpart=0 k2=0 k3=0 k3b=0 w0=2.5u dvt0=1 dvt1=2 dvt2=0 dvt0w=0 dvt1w=0
+  dvt2w=0 dsub=100m minv=50m voffl=0 dvtp0=100p dvtp1=100m lpe0=0 lpeb=0
+  ngate=300e18 nsd=200e18 phin=0 cdsc=0 cdscb=0 cdscd=0 cit=0 voff=-130m
+  etab=0 vfb=-550m u0=49m ua=600p ub=1.2e-18 uc=0 a0=1 ags=0 a1=0 a2=1 b0=0
+  b1=0 keta=40m dwg=0 dwb=0 pclm=20m pdiblc1=1m pdiblc2=1m pdiblcb=-5m
+  drout=500m pvag=10e-21 delta=10m pscbe1=814meg pscbe2=100n fprout=200m
+  pdits=80m pditsd=230m pditsl=2.3meg rsh=5 rsw=80 rdw=80 rdswmin=0 rdwmin=0
+  rswmin=0 prwg=0 prwb=0 wr=1 alpha0=74m alpha1=5m beta0=30 agidl=200u
+  bgidl=2.1g cgidl=200u egidl=800m aigbacc=12m bigbacc=2.8m cigbacc=2m
+  nigbacc=1 aigbinv=14m bigbinv=4m cigbinv=4m eigbinv=1.1 nigbinv=3
+  aigc=15.211m bigc=2.7432m cigc=2m aigsd=15.211m bigsd=2.7432m cigsd=2m
+  nigc=1 poxedge=1 pigcd=1 ntox=1 xrcrg1=12 xrcrg2=5 cgbo=25.6p cgdl=265.3p
+  cgsl=265.3p ckappas=30m ckappad=30m acde=1 moin=15 noff=900m voffcv=20m
+  kt1=-110m kt1l=0 kt2=22m ute=-1.5 ua1=4.31n ub1=7.61e-18 uc1=-56p prt=0
+  at=33k fnoimod=1 tnoimod=0 jss=100u jsws=10p jswgs=100p njs=1 ijthsfwd=10m
+  ijthsrev=1m bvs=10 xjbvs=1 jsd=100u jswd=10p jswgd=100p njd=1 ijthdfwd=10m
+  ijthdrev=1m bvd=10 xjbvd=1 pbs=1 cjs=500u mjs=500m pbsws=1 cjsws=500p
+  mjsws=330m pbswgs=1 cjswgs=300p mjswgs=330m pbd=1 cjd=500u mjd=500m pbswd=1
+  cjswd=500p mjswd=330m pbswgd=1 cjswgd=500p mjswgd=330m tpb=5m tcj=1m
+  tpbsw=5m tcjsw=1m tpbswg=5m tcjswg=1m xtis=3 xtid=3 dmcg=0 dmci=0 dmdg=0
+  dmcgt=0 dwj=0 xgw=0 xgl=0 rshg=400m gbmin=100p rbpb=5 rbpd=15 rbps=15
+  rbdb=15 rbsb=15 ngcon=1
.model PMOS_VTH pmos level=54 version=4.0 binunit=1 paramchk=1 mobmod=0
+  capmod=2 igcmod=1 igbmod=1 geomod=1 diomod=1 rdsmod=0 rbodymod=1 rgatemod=1
+  permod=1 acnqsmod=0 trnqsmod=0 tnom=27 toxe='pToxe' toxp='pToxp' toxm='pToxm' dtox='pdTox'
+  epsrox=3.9 wint=5n lint=3.75n ll=0 wl=0 lln=1 wln=1 lw=0 ww=0 lwn=1 wwn=1
+  lwl=0 wwl=0 xpart=0 toxref='pToxref' vth0=-504.4m k1=400m k2=-10m k3=0 k3b=0
+  w0=2.5u dvt0=1 dvt1=2 dvt2=-32m dvt0w=0 dvt1w=0 dvt2w=0 dsub=100m minv=50m
+  voffl=0 dvtp0=10p dvtp1=50m lpe0=0 lpeb=0 xj=14n ngate=200e18 ndep=2.44e18
+  nsd=200e18 phin=0 cdsc=0 cdscb=0 cdscd=0 cit=0 voff=-126m nfactor=1.8
+  eta0=12.5m etab=0 vfb=550m u0=21m ua=2n ub=500e-21 uc=0 vsat=80k a0=1
+  ags=10e-21 a1=0 a2=1 b0=0 b1=0 keta=-47m dwg=0 dwb=0 pclm=120m pdiblc1=1m
+  pdiblc2=1m pdiblcb=34n drout=560m pvag=10e-21 delta=10m pscbe1=814meg
+  pscbe2=958n fprout=200m pdits=80m pditsd=230m pditsl=2.3meg rsh=5 rdsw=250
+  rsw=75 rdw=75 rdswmin=0 rdwmin=0 rswmin=0 prwg=0 prwb=0 wr=1 alpha0=74m
+  alpha1=5m beta0=30 agidl=200u bgidl=2.1g cgidl=200u egidl=800m aigbacc=12m
+  bigbacc=2.8m cigbacc=2m nigbacc=1 aigbinv=14m bigbinv=4m cigbinv=4m
+  eigbinv=1.1 nigbinv=3 aigc=9.7m bigc=1.25m cigc=800u aigsd=9.7m bigsd=1.25m
+  cigsd=800u nigc=1 poxedge=1 pigcd=1 ntox=1 xrcrg1=12 xrcrg2=5 cgso=110p
+  cgdo=110p cgbo=25.6p cgdl=265.3p cgsl=265.3p ckappas=30m ckappad=30m acde=1
+  moin=15 noff=900m voffcv=20m kt1=-110m kt1l=0 kt2=22m ute=-1.5 ua1=4.31n
+  ub1=7.61e-18 uc1=-56p prt=0 at=33k fnoimod=1 tnoimod=0 jss=100u jsws=10p
+  jswgs=100p njs=1 ijthsfwd=10m ijthsrev=1m bvs=10 xjbvs=1 jsd=100u jswd=10p
+  jswgd=100p njd=1 ijthdfwd=10m ijthdrev=1m bvd=10 xjbvd=1 pbs=1 cjs=500u
+  mjs=500m pbsws=1 cjsws=500p mjsws=330m pbswgs=1 cjswgs=300p mjswgs=330m
+  pbd=1 cjd=500u mjd=500m pbswd=1 cjswd=500p mjswd=330m pbswgd=1 cjswgd=500p
+  mjswgd=330m tpb=5m tcj=1m tpbsw=5m tcjsw=1m tpbswg=5m tcjswg=1m xtis=3
+  xtid=3 dmcg=0 dmci=0 dmdg=0 dmcgt=0 dwj=0 xgw=0 xgl=0 rshg=400m gbmin=100p
+  rbpb=5 rbpd=15 rbps=15 rbdb=15 rbsb=15 ngcon=1
