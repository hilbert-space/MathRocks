.param L = 50n

.param Lnom = 50n
.param Wp = '1.67 * 8 * Lnom'
.param Wn = '8 * Lnom'
.param Lambda = '0.5 * Lnom'

.param Tox = 1n

.param nToxe   = 'Tox + 0.25n'   $ 1.25n
.param nToxp   = 'Tox'           $ 1n
.param nToxm   = 'nToxe'         $ 1.25n
.param nToxref = 'nToxe'         $ 1.25n
.param ndTox   = 'nToxe - nToxp' $ 0.25n

.param pToxe   = 'Tox + 0.3n'    $ 1.3n
.param pToxp   = 'Tox'           $ 1n
.param pToxm   = 'pToxe'         $ 1.3n
.param pToxref = 'pToxe'         $ 1.3n
.param pdTox   = 'pToxe - pToxp' $ 0.3n

.subckt inverter in out dd ss bn bp
M1 out in dd bp pmos
+ L  = 'L'
+ W  = 'Wp'
+ AS = '5 * Wp * Lambda'
+ AD = '5 * Wp * Lambda'
+ PS = '2 * Wp + 10 * Lambda'
+ PD = '2 * Wp + 10 * Lambda'
M2 out in ss bn nmos
+ L  = 'L'
+ W  = 'Wn'
+ AS = '5 * Wn * Lambda'
+ AD = '5 * Wn * Lambda'
+ PS = '2 * Wn + 10 * Lambda'
+ PD = '2 * Wn + 10 * Lambda'
.ends


* PTM High Performance 45nm Metal Gate / High-K / Strained-Si
* nominal Vdd = 1.0V

.model  nmos  nmos  level = 54

+version = 4.0             binunit = 1               paramchk= 1               mobmod  = 0
+capmod  = 2               igcmod  = 1               igbmod  = 1               geomod  = 1
+diomod  = 1               rdsmod  = 0               rbodymod= 1               rgatemod= 1
+permod  = 1               acnqsmod= 0               trnqsmod= 0

+tnom    = 27              toxe    = 'nToxe'         toxp    = 'nToxp'         toxm    = 'nToxm'
+dtox    = 'ndTox'         epsrox  = 3.9             wint    = 5e-009          lint    = 3.75e-009
+ll      = 0               wl      = 0               lln     = 1               wln     = 1
+lw      = 0               ww      = 0               lwn     = 1               wwn     = 1
+lwl     = 0               wwl     = 0               xpart   = 0               toxref  = 'nToxref'
+xl	   = -20e-9

+vth0    = 0.46893         k1      = 0.4             k2      = 0               k3      = 0
+k3b     = 0               w0      = 2.5e-006        dvt0    = 1               dvt1    = 2
+dvt2    = 0               dvt0w   = 0               dvt1w   = 0               dvt2w   = 0
+dsub    = 0.1             minv    = 0.05            voffl   = 0               dvtp0   = 1e-010
+dvtp1   = 0.1             lpe0    = 0               lpeb    = 0               xj      = 1.4e-008
+ngate   = 1e+023          ndep    = 3.24e+018       nsd     = 2e+020          phin    = 0
+cdsc    = 0               cdscb   = 0               cdscd   = 0               cit     = 0
+voff    = -0.13           nfactor = 2.22            eta0    = 0.0055          etab    = 0
+vfb     = -0.55           u0      = 0.054           ua      = 6e-010          ub      = 1.2e-018
+uc      = 0               vsat    = 170000          a0      = 1               ags     = 0
+a1      = 0               a2      = 1               b0      = 0               b1      = 0
+keta    = 0.04            dwg     = 0               dwb     = 0               pclm    = 0.02
+pdiblc1 = 0.001           pdiblc2 = 0.001           pdiblcb = -0.005          drout   = 0.5
+pvag    = 1e-020          delta   = 0.01            pscbe1  = 8.14e+008       pscbe2  = 1e-007
+fprout  = 0.2             pdits   = 0.08            pditsd  = 0.23            pditsl  = 2300000
+rsh     = 5               rdsw    = 155             rsw     = 80              rdw     = 80
+rdswmin = 0               rdwmin  = 0               rswmin  = 0               prwg    = 0
+prwb    = 0               wr      = 1               alpha0  = 0.074           alpha1  = 0.005
+beta0   = 30              agidl   = 0.0002          bgidl   = 2.1e+009        cgidl   = 0.0002
+egidl   = 0.8             aigbacc = 0.012           bigbacc = 0.0028          cigbacc = 0.002
+nigbacc = 1               aigbinv = 0.014           bigbinv = 0.004           cigbinv = 0.004
+eigbinv = 1.1             nigbinv = 3               aigc    = 0.02            bigc    = 0.0025
+cigc    = 0.002           aigsd   = 0.02            bigsd   = 0.0025          cigsd   = 0.002
+nigc    = 1               poxedge = 1               pigcd   = 1               ntox    = 1
+xrcrg1  = 12              xrcrg2  = 5

+cgso    = 1.1e-010        cgdo    = 1.1e-010        cgbo    = 2.56e-011       cgdl    = 2.653e-010
+cgsl    = 2.653e-010      ckappas = 0.03            ckappad = 0.03            acde    = 1
+moin    = 15              noff    = 0.9             voffcv  = 0.02

+kt1     = -0.11           kt1l    = 0               kt2     = 0.022           ute     = -1.5
+ua1     = 4.31e-009       ub1     = 7.61e-018       uc1     = -5.6e-011       prt     = 0
+at      = 33000

+fnoimod = 1               tnoimod = 0

+jss     = 0.0001          jsws    = 1e-011          jswgs   = 1e-010          njs     = 1
+ijthsfwd= 0.01            ijthsrev= 0.001           bvs     = 10              xjbvs   = 1
+jsd     = 0.0001          jswd    = 1e-011          jswgd   = 1e-010          njd     = 1
+ijthdfwd= 0.01            ijthdrev= 0.001           bvd     = 10              xjbvd   = 1
+pbs     = 1               cjs     = 0.0005          mjs     = 0.5             pbsws   = 1
+cjsws   = 5e-010          mjsws   = 0.33            pbswgs  = 1               cjswgs  = 3e-010
+mjswgs  = 0.33            pbd     = 1               cjd     = 0.0005          mjd     = 0.5
+pbswd   = 1               cjswd   = 5e-010          mjswd   = 0.33            pbswgd  = 1
+cjswgd  = 5e-010          mjswgd  = 0.33            tpb     = 0.005           tcj     = 0.001
+tpbsw   = 0.005           tcjsw   = 0.001           tpbswg  = 0.005           tcjswg  = 0.001
+xtis    = 3               xtid    = 3

+dmcg    = 0               dmci    = 0               dmdg    = 0               dmcgt   = 0
+dwj     = 0               xgw     = 0               xgl     = 0

+rshg    = 0.4             gbmin   = 1e-010          rbpb    = 5               rbpd    = 15
+rbps    = 15              rbdb    = 15              rbsb    = 15              ngcon   = 1


.model  pmos  pmos  level = 54

+version = 4.0             binunit = 1               paramchk= 1               mobmod  = 0
+capmod  = 2               igcmod  = 1               igbmod  = 1               geomod  = 1
+diomod  = 1               rdsmod  = 0               rbodymod= 1               rgatemod= 1
+permod  = 1               acnqsmod= 0               trnqsmod= 0

+tnom    = 27              toxe    = 'pToxe'         toxp    = 'pToxp'         toxm    = 'pToxm'
+dtox    = 'pdTox'         epsrox  = 3.9             wint    = 5e-009          lint    = 3.75e-009
+ll      = 0               wl      = 0               lln     = 1               wln     = 1
+lw      = 0               ww      = 0               lwn     = 1               wwn     = 1
+lwl     = 0               wwl     = 0               xpart   = 0               toxref  = 'pToxref'
+xl	   = -20e-9

+vth0    = -0.49158        k1      = 0.4             k2      = -0.01           k3      = 0
+k3b     = 0               w0      = 2.5e-006        dvt0    = 1               dvt1    = 2
+dvt2    = -0.032          dvt0w   = 0               dvt1w   = 0               dvt2w   = 0
+dsub    = 0.1             minv    = 0.05            voffl   = 0               dvtp0   = 1e-011
+dvtp1   = 0.05            lpe0    = 0               lpeb    = 0               xj      = 1.4e-008
+ngate   = 1e+023          ndep    = 2.44e+018       nsd     = 2e+020          phin    = 0
+cdsc    = 0               cdscb   = 0               cdscd   = 0               cit     = 0
+voff    = -0.126          nfactor = 2.1             eta0    = 0.0055          etab    = 0
+vfb     = 0.55            u0      = 0.02            ua      = 2e-009          ub      = 5e-019
+uc      = 0               vsat    = 150000          a0      = 1               ags     = 1e-020
+a1      = 0               a2      = 1               b0      = 0               b1      = 0
+keta    = -0.047          dwg     = 0               dwb     = 0               pclm    = 0.12
+pdiblc1 = 0.001           pdiblc2 = 0.001           pdiblcb = 3.4e-008        drout   = 0.56
+pvag    = 1e-020          delta   = 0.01            pscbe1  = 8.14e+008       pscbe2  = 9.58e-007
+fprout  = 0.2             pdits   = 0.08            pditsd  = 0.23            pditsl  = 2300000
+rsh     = 5               rdsw    = 155             rsw     = 75              rdw     = 75
+rdswmin = 0               rdwmin  = 0               rswmin  = 0               prwg    = 0
+prwb    = 0               wr      = 1               alpha0  = 0.074           alpha1  = 0.005
+beta0   = 30              agidl   = 0.0002          bgidl   = 2.1e+009        cgidl   = 0.0002
+egidl   = 0.8             aigbacc = 0.012           bigbacc = 0.0028          cigbacc = 0.002
+nigbacc = 1               aigbinv = 0.014           bigbinv = 0.004           cigbinv = 0.004
+eigbinv = 1.1             nigbinv = 3               aigc    = 0.010687        bigc    = 0.0012607
+cigc    = 0.0008          aigsd   = 0.010687        bigsd   = 0.0012607       cigsd   = 0.0008
+nigc    = 1               poxedge = 1               pigcd   = 1               ntox    = 1
+xrcrg1  = 12              xrcrg2  = 5

+cgso    = 1.1e-010        cgdo    = 1.1e-010        cgbo    = 2.56e-011       cgdl    = 2.653e-010
+cgsl    = 2.653e-010      ckappas = 0.03            ckappad = 0.03            acde    = 1
+moin    = 15              noff    = 0.9             voffcv  = 0.02

+kt1     = -0.11           kt1l    = 0               kt2     = 0.022           ute     = -1.5
+ua1     = 4.31e-009       ub1     = 7.61e-018       uc1     = -5.6e-011       prt     = 0
+at      = 33000

+fnoimod = 1               tnoimod = 0

+jss     = 0.0001          jsws    = 1e-011          jswgs   = 1e-010          njs     = 1
+ijthsfwd= 0.01            ijthsrev= 0.001           bvs     = 10              xjbvs   = 1
+jsd     = 0.0001          jswd    = 1e-011          jswgd   = 1e-010          njd     = 1
+ijthdfwd= 0.01            ijthdrev= 0.001           bvd     = 10              xjbvd   = 1
+pbs     = 1               cjs     = 0.0005          mjs     = 0.5             pbsws   = 1
+cjsws   = 5e-010          mjsws   = 0.33            pbswgs  = 1               cjswgs  = 3e-010
+mjswgs  = 0.33            pbd     = 1               cjd     = 0.0005          mjd     = 0.5
+pbswd   = 1               cjswd   = 5e-010          mjswd   = 0.33            pbswgd  = 1
+cjswgd  = 5e-010          mjswgd  = 0.33            tpb     = 0.005           tcj     = 0.001
+tpbsw   = 0.005           tcjsw   = 0.001           tpbswg  = 0.005           tcjswg  = 0.001
+xtis    = 3               xtid    = 3

+dmcg    = 0               dmci    = 0               dmdg    = 0               dmcgt   = 0
+dwj     = 0               xgw     = 0               xgl     = 0

+rshg    = 0.4             gbmin   = 1e-010          rbpb    = 5               rbpd    = 15
+rbps    = 15              rbdb    = 15              rbsb    = 15              ngcon   = 1
